`ifndef APB_REGS_PKG__SV
`define APB_REGS_PKG__SV

package apb_regs_pkg;
import uvm_pkg::*;

`include "uvm_macros.svh"

`include "apb_regs.sv"
`include "apb_reg_block.sv"

endpackage : apb_regs_pkg
`endif
