package APB_Package;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "apb_tr.sv"
  `include "apb_cfg.sv"
  `include "apb_seq_list.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_agent.sv"

endpackage : APB_Package
