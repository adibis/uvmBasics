`ifndef APB_TEST_PKG__SV
`define APB_TEST_PKG__SV

package apb_test_pkg;

    import uvm_pkg::*;
    import APB_Package::*;
    import env_pkg::*;


    `include "uvm_macros.svh"

    `include "apb_base_test.sv"
    `include "apb_write_verify_test.sv"
    `include "apb_write_verify_error_test.sv"

endpackage: apb_test_pkg
`endif
