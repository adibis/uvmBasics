`ifndef APB_SEQ_LIST__SV
`define APB_SEQ_LIST__SV

import uvm_pkg::*;

`include "uvm_macros.svh"

`include "apb_base_seq.sv"
`include "apb_read_seq.sv"
`include "apb_write_seq.sv"
`include "apb_write_verify_seq.sv"

`endif
