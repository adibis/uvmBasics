`ifndef APB_REG_PREDICTOR__SV
`define APB_REG_PREDICTOR__SV
typedef uvm_reg_predictor#(apb_seq_item) apb_reg_predictor;
`endif
