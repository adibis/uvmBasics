`ifndef APB_PKG__SV
`define APB_PKG__SV
package apb_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "apb_seq_item.sv"
  `include "apb_cfg.sv"
  `include "apb_seq_list.sv"
  `include "apb_driver.sv"
  `include "apb_monitor.sv"
  `include "apb_reg_adapter.sv"
  `include "apb_reg_predictor.sv"
  `include "apb_agent.sv"

endpackage : apb_pkg
`endif
