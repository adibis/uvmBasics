`ifndef APB_REG_PREDICTOR__SV
`define APB_REG_PREDICTOR__SV
typedef uvm_reg_predictor#(APB_Tr) apb_reg_predictor;
`endif
